magic
tech scmos
timestamp 1524640050
<< checkpaint >>
rect -35 -35 35 35
<< fillm4 >>
rect -5 -5 5 5
<< labels >>
flabel fillm4 0 0 0 0 0 FreeSans 12 0 0 0 PScon
<< end >>
