magic
tech scmos
magscale 1 4
timestamp 1524640050
<< checkpaint >>
rect -114 -130 356 750
use nsubcont  nsubcont_0
timestamp 1524640050
transform 1 0 110 0 1 590
box -40 -40 40 40
use dcont  dcont_0
timestamp 1524640050
transform 1 0 36 0 1 490
box -20 -20 20 20
use dcont  dcont_1
timestamp 1524640050
transform 1 0 36 0 1 450
box -20 -20 20 20
use dcont  dcont_2
timestamp 1524640050
transform 1 0 36 0 1 410
box -20 -20 20 20
use dcont  dcont_3
timestamp 1524640050
transform 1 0 96 0 1 490
box -20 -20 20 20
use dcont  dcont_4
timestamp 1524640050
transform 1 0 96 0 1 450
box -20 -20 20 20
use dcont  dcont_5
timestamp 1524640050
transform 1 0 96 0 1 410
box -20 -20 20 20
use dcont  dcont_6
timestamp 1524640050
transform 1 0 156 0 1 490
box -20 -20 20 20
use dcont  dcont_7
timestamp 1524640050
transform 1 0 156 0 1 450
box -20 -20 20 20
use dcont  dcont_8
timestamp 1524640050
transform 1 0 156 0 1 410
box -20 -20 20 20
use dcont  dcont_9
timestamp 1524640050
transform 1 0 216 0 1 490
box -20 -20 20 20
use dcont  dcont_10
timestamp 1524640050
transform 1 0 216 0 1 450
box -20 -20 20 20
use dcont  dcont_11
timestamp 1524640050
transform 1 0 216 0 1 410
box -20 -20 20 20
use Via  Via_0
timestamp 1524640050
transform 1 0 40 0 1 310
box 0 0 1 1
use pcont  pcont_0
timestamp 1524640050
transform 1 0 40 0 1 310
box -20 -20 20 20
use Via  Via_1
timestamp 1524640050
transform 1 0 220 0 1 260
box 0 0 1 1
use Via  Via_2
timestamp 1524640050
transform 1 0 100 0 1 250
box 0 0 1 1
use pcont  pcont_1
timestamp 1524640050
transform 1 0 100 0 1 250
box -20 -20 20 20
use Via  Via_3
timestamp 1524640050
transform 1 0 160 0 1 180
box 0 0 1 1
use pcont  pcont_2
timestamp 1524640050
transform 1 0 160 0 1 180
box -20 -20 20 20
use dcont  dcont_12
timestamp 1524640050
transform 1 0 36 0 1 74
box -20 -20 20 20
use dcont  dcont_13
timestamp 1524640050
transform 1 0 176 0 1 74
box -20 -20 20 20
use psubcont  psubcont_0
timestamp 1524640050
transform 1 0 100 0 1 10
box -20 -20 20 20
<< labels >>
flabel space 146 198 146 198 2 FreeSans 160 0 0 0 C
flabel space 206 278 206 278 2 FreeSans 160 0 0 0 YB
flabel space 6 20 6 20 2 FreeSans 160 0 0 0 VSS
flabel space 6 570 6 570 2 FreeSans 160 0 0 0 VDD
flabel space 40 328 40 328 2 FreeSans 160 0 0 0 A
flabel space 86 268 86 268 2 FreeSans 160 0 0 0 B
<< end >>
