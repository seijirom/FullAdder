magic
tech scmos
magscale 1 4
timestamp 1524640050
<< checkpaint >>
rect -114 -130 296 750
use nsubcont  nsubcont_0
timestamp 1524640050
transform 1 0 110 0 1 590
box -40 -40 40 40
use dcont  dcont_0
timestamp 1524640050
transform 1 0 46 0 1 490
box -20 -20 20 20
use dcont  dcont_1
timestamp 1524640050
transform 1 0 46 0 1 450
box -20 -20 20 20
use dcont  dcont_2
timestamp 1524640050
transform 1 0 46 0 1 410
box -20 -20 20 20
use dcont  dcont_3
timestamp 1524640050
transform 1 0 146 0 1 490
box -20 -20 20 20
use dcont  dcont_4
timestamp 1524640050
transform 1 0 146 0 1 450
box -20 -20 20 20
use dcont  dcont_5
timestamp 1524640050
transform 1 0 146 0 1 410
box -20 -20 20 20
use Via  Via_0
timestamp 1524640050
transform 1 0 40 0 1 310
box 0 0 1 1
use pcont  pcont_0
timestamp 1524640050
transform 1 0 40 0 1 310
box -20 -20 20 20
use Via  Via_1
timestamp 1524640050
transform 1 0 100 0 1 250
box 0 0 1 1
use pcont  pcont_1
timestamp 1524640050
transform 1 0 100 0 1 250
box -20 -20 20 20
use Via  Via_2
timestamp 1524640050
transform 1 0 160 0 1 190
box 0 0 1 1
use dcont  dcont_6
timestamp 1524640050
transform 1 0 36 0 1 74
box -20 -20 20 20
use dcont  dcont_7
timestamp 1524640050
transform 1 0 96 0 1 74
box -20 -20 20 20
use dcont  dcont_8
timestamp 1524640050
transform 1 0 156 0 1 74
box -20 -20 20 20
use psubcont  psubcont_0
timestamp 1524640050
transform 1 0 100 0 1 10
box -20 -20 20 20
<< labels >>
flabel space 82 266 82 266 2 FreeSans 160 0 0 0 B
flabel space 22 328 22 328 2 FreeSans 160 0 0 0 A
flabel space 6 570 6 570 2 FreeSans 160 0 0 0 VDD
flabel space 6 2 6 2 2 FreeSans 160 0 0 0 VSS
flabel space 148 208 148 208 2 FreeSans 160 0 0 0 YB
<< end >>
