magic
tech scmos
magscale 1 2
timestamp 1521019540
<< checkpaint >>
rect -76 -66 140 270
<< nwell >>
rect -16 96 80 210
<< ntransistor >>
rect 14 12 18 52
rect 24 12 28 52
rect 40 12 44 32
<< ptransistor >>
rect 14 148 18 188
rect 30 148 34 188
rect 46 148 50 188
<< ndiffusion >>
rect 4 51 14 52
rect 12 13 14 51
rect 4 12 14 13
rect 18 12 24 52
rect 28 51 38 52
rect 28 13 30 51
rect 38 13 40 32
rect 28 12 40 13
rect 44 31 54 32
rect 44 13 46 31
rect 44 12 54 13
<< pdiffusion >>
rect 4 187 14 188
rect 12 149 14 187
rect 4 148 14 149
rect 18 187 30 188
rect 18 149 20 187
rect 28 149 30 187
rect 18 148 30 149
rect 34 187 46 188
rect 34 149 36 187
rect 44 149 46 187
rect 34 148 46 149
rect 50 187 60 188
rect 50 149 52 187
rect 50 148 60 149
<< ndcontact >>
rect 4 13 12 51
rect 30 13 38 51
rect 46 13 54 31
<< pdcontact >>
rect 4 149 12 187
rect 20 149 28 187
rect 36 149 44 187
rect 52 149 60 187
<< psubstratepcontact >>
rect -4 -4 4 4
rect 28 -4 36 4
<< nsubstratencontact >>
rect -4 196 4 204
rect 28 196 36 204
<< polysilicon >>
rect 14 188 18 192
rect 30 188 34 192
rect 46 188 50 192
rect 14 82 18 148
rect 30 106 34 148
rect 12 74 18 82
rect 30 78 34 98
rect 14 52 18 74
rect 24 74 34 78
rect 24 52 28 74
rect 46 66 50 148
rect 48 60 50 66
rect 40 32 44 58
rect 14 8 18 12
rect 24 8 28 12
rect 40 8 44 12
<< polycontact >>
rect 26 98 34 106
rect 4 74 12 82
rect 40 58 48 66
<< metal1 >>
rect -4 204 68 206
rect 4 196 28 204
rect 36 196 68 204
rect -4 194 68 196
rect 4 187 12 194
rect 4 148 12 149
rect 20 187 28 188
rect 20 148 28 149
rect 36 187 44 194
rect 36 148 44 149
rect 52 187 60 188
rect 52 148 60 149
rect 22 142 28 148
rect 22 136 46 142
rect 20 106 34 114
rect 4 66 12 74
rect 40 66 46 136
rect 54 134 60 148
rect 52 126 60 134
rect 18 60 40 66
rect 18 58 24 60
rect 6 52 24 58
rect 4 51 12 52
rect 4 12 12 13
rect 30 51 38 52
rect 54 38 60 126
rect 30 6 38 13
rect 46 32 60 38
rect 46 31 54 32
rect 46 12 54 13
rect -4 4 68 6
rect 4 -4 28 4
rect 36 -4 68 4
rect -4 -6 68 -4
<< m1p >>
rect 52 126 60 134
rect 20 106 28 114
rect 4 66 12 74
<< labels >>
rlabel metal1 56 130 56 130 4 Y
rlabel metal1 24 110 24 110 4 B
rlabel metal1 8 200 8 200 4 vdd
rlabel metal1 8 0 8 0 4 gnd
rlabel metal1 8 70 8 70 4 A
<< end >>
