magic
tech scmos
magscale 1 2
timestamp 1521019540
<< checkpaint >>
rect -76 -66 188 270
<< nwell >>
rect -16 96 128 210
<< ntransistor >>
rect 14 12 18 52
rect 32 12 36 32
rect 42 12 46 32
rect 66 12 70 32
rect 76 12 80 32
rect 94 12 98 52
<< ptransistor >>
rect 14 108 18 188
rect 32 148 36 188
rect 42 148 46 188
rect 66 168 70 188
rect 76 168 80 188
rect 94 108 98 188
<< ndiffusion >>
rect 4 51 14 52
rect 12 13 14 51
rect 4 12 14 13
rect 18 51 28 52
rect 18 13 20 51
rect 84 51 94 52
rect 28 13 32 32
rect 18 12 32 13
rect 36 12 42 32
rect 46 30 66 32
rect 46 12 52 30
rect 60 12 66 30
rect 70 12 76 32
rect 80 13 84 32
rect 92 13 94 51
rect 80 12 94 13
rect 98 51 108 52
rect 98 13 100 51
rect 98 12 108 13
<< pdiffusion >>
rect 4 187 14 188
rect 12 109 14 187
rect 4 108 14 109
rect 18 187 32 188
rect 18 109 20 187
rect 28 148 32 187
rect 36 148 42 188
rect 46 187 66 188
rect 46 149 52 187
rect 60 168 66 187
rect 70 168 76 188
rect 80 187 94 188
rect 80 168 84 187
rect 60 149 62 168
rect 46 148 62 149
rect 18 108 28 109
rect 92 109 94 187
rect 84 108 94 109
rect 98 187 108 188
rect 98 109 100 187
rect 98 108 108 109
<< ndcontact >>
rect 4 13 12 51
rect 20 13 28 51
rect 52 12 60 30
rect 84 13 92 51
rect 100 13 108 51
<< pdcontact >>
rect 4 109 12 187
rect 20 109 28 187
rect 52 149 60 187
rect 84 109 92 187
rect 100 109 108 187
<< psubstratepcontact >>
rect -4 -4 4 4
rect 28 -4 36 4
rect 60 -4 68 4
<< nsubstratencontact >>
rect -4 196 4 204
rect 28 196 36 204
rect 60 196 68 204
<< polysilicon >>
rect 14 188 18 192
rect 32 188 36 192
rect 42 188 46 192
rect 66 188 70 192
rect 76 188 80 192
rect 94 188 98 192
rect 14 74 18 108
rect 32 102 36 148
rect 34 96 36 102
rect 30 72 34 94
rect 42 88 46 148
rect 66 146 70 168
rect 62 142 70 146
rect 62 82 66 142
rect 76 114 80 168
rect 30 68 36 72
rect 14 52 18 66
rect 32 32 36 68
rect 42 66 46 80
rect 74 110 80 114
rect 74 84 78 110
rect 42 62 70 66
rect 42 46 44 54
rect 42 32 46 46
rect 66 32 70 62
rect 76 32 80 76
rect 94 52 98 108
rect 14 8 18 12
rect 32 8 36 12
rect 42 8 46 12
rect 66 8 70 12
rect 76 8 80 12
rect 94 8 98 12
<< polycontact >>
rect 26 94 34 102
rect 12 66 20 74
rect 42 80 50 88
rect 58 74 66 82
rect 86 94 94 102
rect 74 76 82 84
rect 44 46 52 54
<< metal1 >>
rect -4 204 116 206
rect 4 196 28 204
rect 36 196 60 204
rect 68 196 116 204
rect -4 194 116 196
rect 4 187 12 188
rect 4 108 12 109
rect 20 187 28 194
rect 50 187 62 188
rect 50 149 52 187
rect 60 149 62 187
rect 50 148 62 149
rect 84 187 92 194
rect 20 108 28 109
rect 36 102 44 114
rect 84 108 92 109
rect 100 187 108 188
rect 4 98 12 100
rect 34 94 44 102
rect 60 94 86 102
rect 12 80 42 86
rect 100 84 108 109
rect 82 76 108 84
rect 20 72 28 74
rect 58 72 66 74
rect 20 66 66 72
rect 44 54 52 66
rect 4 51 12 52
rect 4 12 12 13
rect 20 51 28 52
rect 84 51 92 52
rect 20 6 28 13
rect 50 30 62 32
rect 50 12 52 30
rect 60 12 62 30
rect 84 6 92 13
rect 100 51 108 76
rect 100 12 108 13
rect -4 4 116 6
rect 4 -4 28 4
rect 36 -4 60 4
rect 68 -4 116 4
rect -4 -6 116 -4
<< m2contact >>
rect 52 140 60 148
rect 4 100 12 108
rect 52 94 60 102
rect 4 80 12 88
rect 4 52 12 60
rect 52 32 60 40
<< metal2 >>
rect 4 88 12 100
rect 4 60 12 80
rect 52 102 60 140
rect 52 40 60 94
<< m1p >>
rect 36 106 44 114
rect 100 86 108 94
rect 20 66 28 74
<< labels >>
rlabel metal1 40 110 40 110 4 D
rlabel metal1 104 90 104 90 4 Q
rlabel metal1 8 0 8 0 4 gnd
rlabel metal1 8 200 8 200 4 vdd
rlabel metal1 24 70 24 70 4 CLK
<< end >>
