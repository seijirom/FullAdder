magic
tech scmos
magscale 1 4
timestamp 1524640050
<< checkpaint >>
rect -114 -130 526 750
use nsubcont  nsubcont_0
timestamp 1524640050
transform 1 0 204 0 1 590
box -40 -40 40 40
use dcont  dcont_0
timestamp 1524640050
transform 1 0 36 0 1 516
box -20 -20 20 20
use dcont  dcont_1
timestamp 1524640050
transform 1 0 36 0 1 476
box -20 -20 20 20
use dcont  dcont_2
timestamp 1524640050
transform 1 0 36 0 1 436
box -20 -20 20 20
use dcont  dcont_3
timestamp 1524640050
transform 1 0 96 0 1 516
box -20 -20 20 20
use dcont  dcont_4
timestamp 1524640050
transform 1 0 96 0 1 476
box -20 -20 20 20
use dcont  dcont_5
timestamp 1524640050
transform 1 0 96 0 1 436
box -20 -20 20 20
use dcont  dcont_6
timestamp 1524640050
transform 1 0 156 0 1 516
box -20 -20 20 20
use dcont  dcont_7
timestamp 1524640050
transform 1 0 156 0 1 476
box -20 -20 20 20
use dcont  dcont_8
timestamp 1524640050
transform 1 0 156 0 1 436
box -20 -20 20 20
use dcont  dcont_9
timestamp 1524640050
transform 1 0 226 0 1 516
box -20 -20 20 20
use dcont  dcont_10
timestamp 1524640050
transform 1 0 226 0 1 476
box -20 -20 20 20
use dcont  dcont_11
timestamp 1524640050
transform 1 0 226 0 1 436
box -20 -20 20 20
use dcont  dcont_12
timestamp 1524640050
transform 1 0 326 0 1 516
box -20 -20 20 20
use dcont  dcont_13
timestamp 1524640050
transform 1 0 326 0 1 476
box -20 -20 20 20
use dcont  dcont_14
timestamp 1524640050
transform 1 0 326 0 1 436
box -20 -20 20 20
use dcont  dcont_15
timestamp 1524640050
transform 1 0 386 0 1 516
box -20 -20 20 20
use dcont  dcont_16
timestamp 1524640050
transform 1 0 386 0 1 476
box -20 -20 20 20
use dcont  dcont_17
timestamp 1524640050
transform 1 0 386 0 1 436
box -20 -20 20 20
use Via  Via_0
timestamp 1524640050
transform 1 0 140 0 1 294
box 0 0 1 1
use pcont  pcont_0
timestamp 1524640050
transform 1 0 140 0 1 294
box -20 -20 20 20
use pcont  pcont_1
timestamp 1524640050
transform 1 0 286 0 1 294
box -20 -20 20 20
use Via  Via_1
timestamp 1524640050
transform 1 0 390 0 1 270
box 0 0 1 1
use Via  Via_2
timestamp 1524640050
transform 1 0 80 0 1 234
box 0 0 1 1
use pcont  pcont_2
timestamp 1524640050
transform 1 0 80 0 1 234
box -20 -20 20 20
use pcont  pcont_3
timestamp 1524640050
transform 1 0 226 0 1 234
box -20 -20 20 20
use pcont  pcont_4
timestamp 1524640050
transform 1 0 346 0 1 174
box -20 -20 20 20
use dcont  dcont_18
timestamp 1524640050
transform 1 0 36 0 1 74
box -20 -20 20 20
use dcont  dcont_19
timestamp 1524640050
transform 1 0 136 0 1 74
box -20 -20 20 20
use dcont  dcont_20
timestamp 1524640050
transform 1 0 206 0 1 74
box -20 -20 20 20
use dcont  dcont_21
timestamp 1524640050
transform 1 0 266 0 1 74
box -20 -20 20 20
use dcont  dcont_22
timestamp 1524640050
transform 1 0 326 0 1 74
box -20 -20 20 20
use dcont  dcont_23
timestamp 1524640050
transform 1 0 386 0 1 74
box -20 -20 20 20
use psubcont  psubcont_0
timestamp 1524640050
transform 1 0 204 0 1 10
box -20 -20 20 20
<< labels >>
flabel space 140 288 140 288 2 FreeSans 160 0 0 0 A
flabel space 80 228 80 228 2 FreeSans 160 0 0 0 B
flabel space 6 570 6 570 2 FreeSans 160 0 0 0 VDD
flabel space 6 20 6 20 2 FreeSans 160 0 0 0 VSS
flabel space 380 282 380 282 2 FreeSans 160 0 0 0 YB
<< end >>
