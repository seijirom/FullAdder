magic
tech scmos
magscale 1 4
timestamp 1524640050
<< checkpaint >>
rect -114 -130 656 750
use nsubcont  nsubcont_0
timestamp 1524640050
transform 1 0 100 0 1 590
box -40 -40 40 40
use nsubcont  nsubcont_1
timestamp 1524640050
transform 1 0 382 0 1 590
box -40 -40 40 40
use dcont  dcont_0
timestamp 1524640050
transform 1 0 36 0 1 490
box -20 -20 20 20
use dcont  dcont_1
timestamp 1524640050
transform 1 0 36 0 1 450
box -20 -20 20 20
use dcont  dcont_2
timestamp 1524640050
transform 1 0 36 0 1 410
box -20 -20 20 20
use dcont  dcont_3
timestamp 1524640050
transform 1 0 96 0 1 490
box -20 -20 20 20
use dcont  dcont_4
timestamp 1524640050
transform 1 0 96 0 1 450
box -20 -20 20 20
use dcont  dcont_5
timestamp 1524640050
transform 1 0 96 0 1 410
box -20 -20 20 20
use dcont  dcont_6
timestamp 1524640050
transform 1 0 156 0 1 490
box -20 -20 20 20
use dcont  dcont_7
timestamp 1524640050
transform 1 0 156 0 1 450
box -20 -20 20 20
use dcont  dcont_8
timestamp 1524640050
transform 1 0 156 0 1 410
box -20 -20 20 20
use dcont  dcont_9
timestamp 1524640050
transform 1 0 216 0 1 490
box -20 -20 20 20
use dcont  dcont_10
timestamp 1524640050
transform 1 0 216 0 1 450
box -20 -20 20 20
use dcont  dcont_11
timestamp 1524640050
transform 1 0 216 0 1 410
box -20 -20 20 20
use dcont  dcont_12
timestamp 1524640050
transform 1 0 276 0 1 490
box -20 -20 20 20
use dcont  dcont_13
timestamp 1524640050
transform 1 0 276 0 1 450
box -20 -20 20 20
use dcont  dcont_14
timestamp 1524640050
transform 1 0 276 0 1 410
box -20 -20 20 20
use dcont  dcont_15
timestamp 1524640050
transform 1 0 336 0 1 490
box -20 -20 20 20
use dcont  dcont_16
timestamp 1524640050
transform 1 0 336 0 1 450
box -20 -20 20 20
use dcont  dcont_17
timestamp 1524640050
transform 1 0 336 0 1 410
box -20 -20 20 20
use dcont  dcont_18
timestamp 1524640050
transform 1 0 396 0 1 490
box -20 -20 20 20
use dcont  dcont_19
timestamp 1524640050
transform 1 0 396 0 1 450
box -20 -20 20 20
use dcont  dcont_20
timestamp 1524640050
transform 1 0 396 0 1 410
box -20 -20 20 20
use dcont  dcont_21
timestamp 1524640050
transform 1 0 456 0 1 490
box -20 -20 20 20
use dcont  dcont_22
timestamp 1524640050
transform 1 0 456 0 1 450
box -20 -20 20 20
use dcont  dcont_23
timestamp 1524640050
transform 1 0 456 0 1 410
box -20 -20 20 20
use dcont  dcont_24
timestamp 1524640050
transform 1 0 516 0 1 490
box -20 -20 20 20
use dcont  dcont_25
timestamp 1524640050
transform 1 0 516 0 1 450
box -20 -20 20 20
use dcont  dcont_26
timestamp 1524640050
transform 1 0 516 0 1 410
box -20 -20 20 20
use Via  Via_0
timestamp 1524640050
transform 1 0 40 0 1 310
box 0 0 1 1
use pcont  pcont_0
timestamp 1524640050
transform 1 0 40 0 1 310
box -20 -20 20 20
use Via  Via_1
timestamp 1524640050
transform 1 0 460 0 1 230
box 0 0 1 1
use dcont  dcont_27
timestamp 1524640050
transform 1 0 36 0 1 74
box -20 -20 20 20
use dcont  dcont_28
timestamp 1524640050
transform 1 0 96 0 1 74
box -20 -20 20 20
use dcont  dcont_29
timestamp 1524640050
transform 1 0 156 0 1 74
box -20 -20 20 20
use dcont  dcont_30
timestamp 1524640050
transform 1 0 216 0 1 74
box -20 -20 20 20
use dcont  dcont_31
timestamp 1524640050
transform 1 0 276 0 1 74
box -20 -20 20 20
use dcont  dcont_32
timestamp 1524640050
transform 1 0 336 0 1 74
box -20 -20 20 20
use dcont  dcont_33
timestamp 1524640050
transform 1 0 396 0 1 74
box -20 -20 20 20
use dcont  dcont_34
timestamp 1524640050
transform 1 0 456 0 1 74
box -20 -20 20 20
use dcont  dcont_35
timestamp 1524640050
transform 1 0 516 0 1 74
box -20 -20 20 20
use psubcont  psubcont_0
timestamp 1524640050
transform 1 0 100 0 1 10
box -20 -20 20 20
use psubcont  psubcont_1
timestamp 1524640050
transform 1 0 366 0 1 10
box -20 -20 20 20
<< labels >>
flabel space 452 248 452 248 2 FreeSans 160 0 0 0 YB
flabel space 6 20 6 20 2 FreeSans 160 0 0 0 VSS
flabel space 6 570 6 570 2 FreeSans 160 0 0 0 VDD
flabel space 40 328 40 328 2 FreeSans 160 0 0 0 A
<< end >>
