magic
tech scmos
magscale 1 4
timestamp 1524640050
<< checkpaint >>
rect -114 -130 356 750
use nsubcont  nsubcont_0
timestamp 1524640050
transform 1 0 164 0 1 590
box -40 -40 40 40
use dcont  dcont_0
timestamp 1524640050
transform 1 0 56 0 1 490
box -20 -20 20 20
use dcont  dcont_1
timestamp 1524640050
transform 1 0 56 0 1 450
box -20 -20 20 20
use dcont  dcont_2
timestamp 1524640050
transform 1 0 56 0 1 410
box -20 -20 20 20
use dcont  dcont_3
timestamp 1524640050
transform 1 0 156 0 1 490
box -20 -20 20 20
use dcont  dcont_4
timestamp 1524640050
transform 1 0 156 0 1 450
box -20 -20 20 20
use dcont  dcont_5
timestamp 1524640050
transform 1 0 156 0 1 410
box -20 -20 20 20
use dcont  dcont_6
timestamp 1524640050
transform 1 0 216 0 1 490
box -20 -20 20 20
use dcont  dcont_7
timestamp 1524640050
transform 1 0 216 0 1 450
box -20 -20 20 20
use dcont  dcont_8
timestamp 1524640050
transform 1 0 216 0 1 410
box -20 -20 20 20
use Via  Via_0
timestamp 1524640050
transform 1 0 40 0 1 310
box 0 0 1 1
use pcont  pcont_0
timestamp 1524640050
transform 1 0 40 0 1 310
box -20 -20 20 20
use Via  Via_1
timestamp 1524640050
transform 1 0 100 0 1 250
box 0 0 1 1
use pcont  pcont_1
timestamp 1524640050
transform 1 0 100 0 1 250
box -20 -20 20 20
use Via  Via_2
timestamp 1524640050
transform 1 0 160 0 1 260
box 0 0 1 1
use pcont  pcont_2
timestamp 1524640050
transform 1 0 160 0 1 260
box -20 -20 20 20
use Via  Via_3
timestamp 1524640050
transform 1 0 220 0 1 190
box 0 0 1 1
use dcont  dcont_9
timestamp 1524640050
transform 1 0 36 0 1 110
box -20 -20 20 20
use dcont  dcont_10
timestamp 1524640050
transform 1 0 96 0 1 110
box -20 -20 20 20
use dcont  dcont_11
timestamp 1524640050
transform 1 0 156 0 1 110
box -20 -20 20 20
use dcont  dcont_12
timestamp 1524640050
transform 1 0 216 0 1 110
box -20 -20 20 20
use psubcont  psubcont_0
timestamp 1524640050
transform 1 0 130 0 1 10
box -20 -20 20 20
<< labels >>
flabel space 202 208 202 208 2 FreeSans 160 0 0 0 YB
flabel space 160 254 160 254 2 FreeSans 160 0 0 0 B0
flabel space 6 20 6 20 2 FreeSans 160 0 0 0 VSS
flabel space 6 570 6 570 2 FreeSans 160 0 0 0 VDD
flabel space 40 304 40 304 2 FreeSans 160 0 0 0 A0
flabel space 100 244 100 244 2 FreeSans 160 0 0 0 A1
<< end >>
